module tb;
  initial begin
    repeat(5) begin
      $display("Hello World!");
    end
  end
endmodule
